
--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY PROGRAM_COUNTER IS
	PORT (D : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			Q : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			RESET : IN STD_LOGIC;
			CLK : IN STD_LOGIC);
END PROGRAM_COUNTER; 



ARCHITECTURE BEHAVIORAL OF PROGRAM_COUNTER IS

SIGNAL Q_INT: STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');

BEGIN

PROCESS(CLK,RESET,D)
BEGIN

		IF RESET = '1' THEN
		Q_INT <= (OTHERS => '0');  --ASYNCRONOUS INPUT CLEARS THE VECTOR
		ELSIF FALLING_EDGE(CLK) THEN
		Q_INT <= D;
		ELSE 
			NULL;
		END IF;
END PROCESS;
Q <= Q_INT;   							--CONCURRENT STATEMENT

END BEHAVIORAL;

