--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
LIBRARY IEEE;


USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ROM_MEMORY IS
PORT ( ADDRESS : IN STD_LOGIC_VECTOR ( 4 DOWNTO 0 );  --ALLOCATE 32 REGISTERS
		 DATA : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 0 ));  --2 BYTE DATA
END ROM_MEMORY;

ARCHITECTURE BEHAVIORAL OF ROM_MEMORY IS
BEGIN

PROCESS(ADDRESS)

SUBTYPE ROM_REGISTER IS STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
TYPE ROM_WIDTH IS ARRAY ( 0 TO 31 ) OF ROM_REGISTER;
VARIABLE ROM : ROM_WIDTH := ( "0001000100010001" , "1010101010101010" , "1000111011101010" , "0010101010101010" , "0000101010101010" ,OTHERS => ( OTHERS => '0' ) );

VARIABLE ADDRESS_INT : NATURAL;

BEGIN

ADDRESS_INT := TO_INTEGER(UNSIGNED(ADDRESS));
DATA <= ROM(ADDRESS_INT);

END PROCESS;
END BEHAVIORAL;



