--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY MUX_2X1 IS
	PORT (E: IN STD_LOGIC; 
			DATA1 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);  --Datos]
			DATA2 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			DATA_OUT: OUT STD_LOGIC_VECTOR (31 DOWNTO 0));		
END MUX_2X1; 

ARCHITECTURE BEHAVIORAL OF MUX_2X1 IS

BEGIN
DATA_OUT <= DATA1 WHEN E= '1' ELSE DATA2;
		
END BEHAVIORAL;

