--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ALU IS
	PORT (CTL: IN STD_LOGIC_VECTOR(2 DOWNTO 0); 
			A : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			B : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ZERO : OUT STD_LOGIC;
			RESULT: OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
			
END ALU; 

ARCHITECTURE BEHAVIORAL OF ALU IS
	SIGNAL sRESULT : UNSIGNED (31 DOWNTO 0) := (OTHERS => '0');
BEGIN

PROCESS(A,B,CTL)
BEGIN

	CASE CTL IS 
		WHEN "000" => sRESULT <= UNSIGNED(A AND B); --A & B
		WHEN "001" => sRESULT <= UNSIGNED(A OR B);  --A || B
		WHEN "010" => sRESULT <= UNSIGNED(SIGNED(A) + SIGNED(B));
		WHEN "011" => sRESULT <= UNSIGNED(A);
		WHEN "100" => sRESULT <= UNSIGNED(B(15 DOWNTO 0)) & x"0000";
		WHEN "101" => NULL;
		WHEN "110" => sRESULT <= UNSIGNED(SIGNED(A) - SIGNED(B));
		WHEN "111" => 
		
							IF (A < B) THEN
								sRESULT <= x"00000001";
								
							ELSE
								sRESULT <= (OTHERS => '0');
							END IF;
		  	
	END CASE;
END PROCESS;


   ZERO <= '1' WHEN sRESULT = x"00000000" ELSE '0';

	RESULT <= STD_LOGIC_VECTOR(sRESULT);
	
END BEHAVIORAL;
		
