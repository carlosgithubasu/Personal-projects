LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY VGA IS
	PORT (
		CLK50M    : IN STD_LOGIC;
		RESET		 : IN STD_LOGIC;
		VIDEO_ON  : OUT STD_LOGIC;
		COLUMN    : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		ROW       : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		HS        : OUT STD_LOGIC;
		VS        : OUT STD_LOGIC
	);
END VGA;

ARCHITECTURE BEHAVIORAL OF VGA IS

	-- HORIZONTAL SYNC PARAMETERS:
	
	CONSTANT TS_H : INTEGER := 800;
	CONSTANT TDISP_H : INTEGER := 640;
	CONSTANT TPW_H : INTEGER := 96;
	CONSTANT TFP_H : INTEGER := 16;
	CONSTANT TBP_H : INTEGER := 48;
	

	-- VERTICAL SYNC PARAMETERS:
	
	CONSTANT TS_V : INTEGER := 521;
	CONSTANT TDISP_V : INTEGER := 480;
	CONSTANT TPW_V : INTEGER := 2;
	CONSTANT TFP_V : INTEGER := 10;
	CONSTANT TBP_V : INTEGER := 29;

	-- SIGNALS AND COUNTERS:

	SIGNAL CLK25M : STD_LOGIC := '0';
	SIGNAL COUNTER_H : INTEGER RANGE 0 TO 799 := 0;
	SIGNAL NEXT_COUNTER_H : INTEGER RANGE 0 TO 799 := 0;
	SIGNAL COUNTER_V : INTEGER RANGE 0 TO 520 := 0;

BEGIN
	PROCESS (CLK50M)
	BEGIN
		IF (RISING_EDGE(CLK50M)) THEN
			CLK25M <= NOT CLK25M;
		END IF;
	END PROCESS;

	PROCESS (CLK25M, RESET)
	BEGIN
		IF RESET = '1' THEN
			COUNTER_H <= 0;
		ELSIF (RISING_EDGE(CLK25M)) THEN
			COUNTER_H <= NEXT_COUNTER_H;
		END IF;
	END PROCESS;

	NEXT_COUNTER_H <= (COUNTER_H + 1) WHEN (COUNTER_H < TS_H - 1) ELSE 0;

	PROCESS (CLK25M, RESET)
	BEGIN
		IF RESET = '1' THEN
			COUNTER_V <= 0;
		ELSIF (RISING_EDGE(CLK25M)) THEN
			IF (NEXT_COUNTER_H = 0) THEN
				IF (COUNTER_V = TS_V - 1) THEN
					COUNTER_V <= 0;
				ELSE
					COUNTER_V <= COUNTER_V + 1;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	HS <= '0' WHEN (COUNTER_H < TPW_H) ELSE '1';
	VS <= '0' WHEN (COUNTER_V < TPW_V) ELSE '1';

	VIDEO_ON <= '0' WHEN ((COUNTER_H < TPW_H + TBP_H) OR (COUNTER_H > TDISP_H + TPW_H + TBP_H - 1 ) OR (COUNTER_V < TPW_V + TBP_V) OR (COUNTER_V > TDISP_V + TPW_V + TBP_V - 1)) ELSE '1';
	
	COLUMN <= CONV_STD_LOGIC_VECTOR(COUNTER_H,10);
	ROW <= CONV_STD_LOGIC_VECTOR(COUNTER_V,10);
	
	
END BEHAVIORAL;