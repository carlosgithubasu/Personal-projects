--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY DATA_MEMORY IS
	PORT( ADDRESS : IN STD_LOGIC_VECTOR (4 DOWNTO 0 );
			WRITE_DATA : IN STD_LOGIC_VECTOR (31 DOWNTO 0 );
			READ_DATA : OUT STD_LOGIC_VECTOR (31 DOWNTO 0 );
			CLK, WRITE_ENABLE, READ_ENABLE, ENABLE: IN STD_LOGIC);
END  DATA_MEMORY;

ARCHITECTURE BEHAVIORAL OF DATA_MEMORY IS

SUBTYPE DATA_MEMORY_REGISTER IS STD_LOGIC_VECTOR ( 31 DOWNTO 0 );      --Ancho del bus memoria de datos
TYPE DATA_MEMORY_WIDTH IS ARRAY ( 0 TO 31 ) OF  DATA_MEMORY_REGISTER;  --Ancho del bus de direcciones
SIGNAL MEMORY_DATA : DATA_MEMORY_WIDTH := ( OTHERS => (OTHERS => '0'));--relleno direcciones con 0'S

SIGNAL RD : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');


BEGIN

PROCESS(CLK, WRITE_ENABLE,READ_ENABLE)
BEGIN

  IF FALLING_EDGE(CLK) THEN
		
		IF WRITE_ENABLE  = '1' AND READ_ENABLE = '0' THEN
		MEMORY_DATA (TO_INTEGER(UNSIGNED(ADDRESS(6 DOWNTO 2)))) <=  WRITE_DATA;
		RD <= (OTHERS => '0');
		ELSIF WRITE_ENABLE = '0' AND READ_ENABLE = '1' THEN
		RD <= MEMORY_DATA (TO_INTEGER(UNSIGNED(ADDRESS(6 DOWNTO 2))));
		ELSE
				RD <= (OTHERS => '0');
		END IF;
  END IF;
END PROCESS;


	READ_DATA <= RD;
	
END BEHAVIORAL;
		
