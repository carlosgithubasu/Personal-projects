

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY lcd_controller IS
	PORT (
		clk : IN STD_LOGIC; 
		reset_n : IN STD_LOGIC; 
		lcd_enable : IN STD_LOGIC; 
		lcd_bus : IN STD_LOGIC_VECTOR(9 DOWNTO 0); 
		busy : OUT STD_LOGIC := '1'; 
		rw, rs, e : OUT STD_LOGIC; 
		lcd_data : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
	
	
END lcd_controller;

ARCHITECTURE controller OF lcd_controller IS
	TYPE CONTROL IS(power_up, initialize, ready, send);
	SIGNAL state : CONTROL;
	CONSTANT freq : INTEGER := 50;
BEGIN
	PROCESS (clk)
VARIABLE clk_count : INTEGER := 0;
BEGIN
	IF (clk'EVENT AND clk = '1') THEN
 

		CASE state IS
 
 
			WHEN power_up => 
				busy <= '1';
				IF (clk_count < (50000 * freq)) THEN --wait 50 ms
					clk_count := clk_count + 1;
					state <= power_up;
				ELSE --power-up complete
					clk_count := 0;
					rs <= '0';
					rw <= '0';
					lcd_data <= "00110000";
					state <= initialize;
				END IF;
 
				--cycle through initialization sequence 
			WHEN initialize => 
				busy <= '1';
				clk_count := clk_count + 1;
				IF (clk_count < (10 * freq)) THEN --function set   wait 10 us
					lcd_data <= "00111100"; --2-line mode, display on
 
					e <= '1';
					state <= initialize;
				ELSIF (clk_count < (60 * freq)) THEN --wait 50 us
					lcd_data <= "00000000";
					e <= '0';
					state <= initialize;
				ELSIF (clk_count < (70 * freq)) THEN --display on/off control 10 us
					lcd_data <= "00001100"; --display on, cursor off, blink off
 
					e <= '1';
					state <= initialize;
				ELSIF (clk_count < (120 * freq)) THEN --wait 50 us
					lcd_data <= "00000000";
					e <= '0';
					state <= initialize;   ; -- 10us
				ELSIF (clk_count < (130 * freq)) THEN --display clear
					lcd_data <= "00000001";
					e <= '1';
					state <= initialize;
				ELSIF (clk_count < (2130 * freq)) THEN --wait 2 ms
					lcd_data <= "00000000";
					e <= '0';
					state <= initialize;
				ELSIF (clk_count < (2140 * freq)) THEN --entry mode set
					lcd_data <= "00000110"; --increment mode, entire shift off
 
					e <= '1';
					state <= initialize;
				ELSIF (clk_count < (2200 * freq)) THEN --wait 60 us
					lcd_data <= "00000000";
					e <= '0';
					state <= initialize;
				ELSE --initialization complete
					clk_count := 0;
					busy <= '0'; 
					state <= ready;
				END IF; 
 
				--wait for the enable signal and then latch in the instruction
			WHEN ready => 
				IF (lcd_enable = '1') THEN
					busy <= '1';
					rs <= lcd_bus(9);
					rw <= lcd_bus(8);
					lcd_data <= lcd_bus(7 DOWNTO 0);
					clk_count := 0; 
					state <= send;
				ELSE
					busy <= '0';
					rs <= '0';
					rw <= '0';
					lcd_data <= "00000000";
					clk_count := 0;
					state <= ready;
				END IF;
 
				--send instruction to lcd 
			WHEN send => 
				busy <= '1';
				IF (clk_count < (50 * freq)) THEN --do not exit for 50us
					busy <= '1';
					IF (clk_count < freq) THEN --negative enable
						e <= '0';
					ELSIF (clk_count < (14 * freq)) THEN --positive enable half-cycle
						e <= '1';
					ELSIF (clk_count < (27 * freq)) THEN --negative enable half-cycle
						e <= '0';
					END IF;
					clk_count := clk_count + 1;
					state <= send;
				ELSE
					clk_count := 0;
					state <= ready;
				END IF;

		END CASE; 
 
		--reset
		IF (reset_n = '0') THEN
			state <= power_up;
		END IF;
 
	END IF;
END PROCESS;
END controller;