--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ADD IS 
PORT( A,B : IN STD_LOGIC_VECTOR ( 31 DOWNTO 0);  -- DATA INPUTS A & B
		C : OUT STD_LOGIC_VECTOR ( 31 DOWNTO 0);   -- 31 DOWN TO 0 => OVERFLOW ?
      CARRY_OUT : OUT STD_LOGIC);                --CARRY OUT
		END ADD;

ARCHITECTURE EQUATIONS OF ADD IS

BEGIN
		C  <=  STD_LOGIC_VECTOR(UNSIGNED(A) + UNSIGNED(B));
END EQUATIONS;



   