
--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
--DONE
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY SIGN_EXTENDER IS
	PORT (A: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			B : OUT STD_LOGIC_VECTOR (31 DOWNTO 0));
END SIGN_EXTENDER; 

ARCHITECTURE BEHAVIORAL OF SIGN_EXTENDER IS

BEGIN
    B <= (31 DOWNTO 16 => A(15)) & A;
END BEHAVIORAL;

