LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DEBOUNCEDEVOLUTION IS
	PORT (
		CLK   : IN STD_LOGIC;
		DIN   : IN STD_LOGIC;
		QOUT  : OUT STD_LOGIC
	);
END DEBOUNCEDEVOLUTION;

ARCHITECTURE Behavioral OF DEBOUNCEDEVOLUTION IS
	SIGNAL Q1, Q2, Q3 : STD_LOGIC;
BEGIN
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			Q1 <= DIN;
			Q2 <= Q1;
			Q3 <= Q2;
		END IF;
	END PROCESS;

	QOUT <= Q1 AND Q2 AND  Q3;

END Behavioral;