LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY CLK1KHZ IS
	PORT (
		MCLK : IN STD_LOGIC;
		CLKOUT : OUT STD_LOGIC
	);
END CLK1KHZ;

ARCHITECTURE Behavioral OF CLK1KHZ IS
	
SIGNAL CLK1KHZ : STD_LOGIC:='0';
	
BEGIN
	PROCESS (MCLK)
	VARIABLE COUNTER : INTEGER := 0;
	BEGIN
		IF MCLK = '1' AND MCLK'EVENT THEN
			IF COUNTER = 25000 THEN
				COUNTER := 0;
				CLK1KHZ <= NOT CLK1KHZ;
			ELSE COUNTER := COUNTER + 1;
			END IF;
		ELSE NULL;
		END IF;
	END PROCESS;

	CLKOUT <= CLK1KHZ;
END Behavioral;