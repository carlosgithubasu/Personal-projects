--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;


ENTITY RAM_MEMORY IS 
	PORT( ADDRESS : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0 );       --ALLOCATE 16 REGISTERS
			WRITE_DATA : IN STD_LOGIC_VECTOR ( 15 DOWNTO 0 );   --2 BYTE DATA
			READ_DATA : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 0 );
			RW , CLK : IN  STD_LOGIC);                          --READ/WRITE AND CLOCK SIGNAL
END RAM_MEMORY;


ARCHITECTURE BEHAVIORAL OF  RAM_MEMORY IS

SUBTYPE RAM_REGISTER IS STD_LOGIC_VECTOR ( 15 DOWNTO 0 );  --DATA BUS WIDTH
TYPE REG_WIDTH IS ARRAY ( 0 TO 15 ) OF  RAM_REGISTER;  	  --16 ALLOCATIONS
SIGNAL  RAM : REG_WIDTH := ( OTHERS => (OTHERS => '0')); 

SIGNAL RD : STD_LOGIC_VECTOR(15 DOWNTO 0):= (OTHERS =>'0'); --SIGNAL WHAT FOR?

BEGIN 
PROCESS(CLK,RW)   
			  
BEGIN

	IF RISING_EDGE(CLK) THEN
		IF RW = '0'  THEN
		RAM ( TO_INTEGER(  UNSIGNED( ADDRESS) ) ) <= WRITE_DATA;  --WRITE RAM WHEN '0'
		ELSIF RW = '1' THEN
	   
		READ_DATA <= RAM( TO_INTEGER ( UNSIGNED (ADDRESS) ) );    --READ FROM RAM WHEN  '1'
		
		ELSE NULL;  
		
		END IF;
	END IF;
END PROCESS;

READ_DATA <= RD;

END BEHAVIORAL;

		
		
	


