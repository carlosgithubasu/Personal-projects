--Carlos Perez Araujo , Tecnologico de Estudios Superiores de Monterrey
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY TEST_keypad IS
END TEST_keypad;

ARCHITECTURE TEST OF TEST_keypad IS

	COMPONENT TESTING_KEYPAD IS
	PORT (
		CLK : IN STD_LOGIC;
		ROW : IN STD_LOGIC_VECTOR(0 TO 3);
		COL : OUT STD_LOGIC_VECTOR(0 TO 3);
	   KEY : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	   KEY_AVAILABLE : OUT STD_LOGIC
		
	);
END COMPONENT;
	
	
SIGNAL CLK : STD_LOGIC;
SIGNAL ROW : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL COL : STD_LOGIC_VECTOR(0 TO 3);
SIGNAL KEY : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL KEY_AVAILABLE :  STD_LOGIC;

	
	
BEGIN
	PORTMAP : TESTING_KEYPAD
	PORT MAP ( CLK => CLK , ROW => ROW, COL => COL , KEY => KEY , KEY_AVAILABLE => KEY_AVAILABLE);

STIMULUS : 
PROCESS
BEGIN
	clk <= '0';
	WAIT FOR 10 ns;

	clk <= '1';
	ROW <= "0001";
	

	WAIT FOR 10 ns;
	clk <= '0';
	WAIT FOR 10 ns;
	clk <= '1';

	WAIT FOR 10 ns;
	clk <= '0';
	

	WAIT FOR 10 ns;
	clk <= '1';
	
	WAIT FOR 10 ns;
	clk <= '0';
	ROW <= "0100";

END PROCESS;
END TEST;
