library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;

--VHDL CODE FOR 4BIT ADDER USING THE STD_LOGICC_UNSIGNED PACKAGE

entity Adder_4 is 
	port(A,B: IN STD_LOGIC_VECTOR(3 DOWNTO 0); CI: IN STD_LOGIC; --INPUTS
		S:OUT STD_LOGIC_VECTOR(3 DOWNTO 0); CO: OUT STD_LOGIC);
END ADDER_4;

ARCHITECTURE OVERLOAD OF ADDER_4 IS
SIGNAL SUM5 : STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN

SUM5 <= '0' & A + B + CI; --ADDER
S<= SUM5(3 DOWNTO 0);
CO<= SUM5(4);
END OVERLOAD;